// RAM Model
//
// +-----------------------------+
// |    Copyright 1996 DOULOS    |
// |       Library: Memory       |
// |   designer : John Aynsley   |
// +-----------------------------+

module RamChip (Address, Data, CS, WE, OE);

parameter AddressSize = 1;
parameter WordSize = 1;

input [AddressSize-1:0] Address;
inout [WordSize-1:0] Data;
input CS, WE, OE;

reg [WordSize-1:0] Mem [0:1<<AddressSize];

assign Data = (!CS && !OE) ? Mem[Address] : {WordSize{1'bz}};

always @(CS or WE)
  if (!CS && !WE)
    Mem[Address] = Data;

always @(WE or OE)
  if (!WE && !OE)
    $display("Operational error in RamChip: OE and WE both active");

endmodule // RamChip



interface ramIff (input clk);

   logic 	   CS, WE, OE;
   logic [3:0] 	   Address;
   logic [7:0] 	   Data;

   clocking cb @(posedge clk);
      input 	   Data;
      output 	   CS, WE, OE, Address;
      
endclocking
 	   

endinterface // ramIff

class driver;
   virtual     ramIff vif;
   Packet pkt;
   Packet pkt_q[$];
   
   function new(ramIff vif);
      this.vif = vif;
      
   endfunction // new
   
   task send_rqt(input pkt);
      pkt_q.push_back(pkt);
      
      vif.cb.CS <= pkt.CS;
      vif.cb.WE <= pkt.WE;
      vif.cb.OE <= pkt.OE;
      vif.cb.Address <= pkt.Address;
      vif.cb.Data <= pkt.Data;
      @vif.cb;
      
   endtask // send_rqt
endclass // driver

class oMonitor;
   virtual ramIff vif;
   logic [7:0] Data_q[$];
   
   function new();
      fork
	 captureOp();
      join_none
      
   endfunction // new
      
   task captureOp ()  ;
      if(vif.cb.WE)begin
	 @vif.cb;
	 #1
	 Data_q.push_back(vif.Data);
      end
      
   endtask // captureOp
   
endclass // oMonitor

class Packet;
//Create randomized packet.

   rand logic CS, WE, OE;
   rand logic [7:0] Data;
   rand logic [4:0] Address;

   constraint configCon {
      CS == 1;
      if(WE==1)(OE==0);
   }

   
endclass // Packet




module top;

   logic clock;

   //Interface
   ramIff iftest(clk);
   //Components
   oMonitor mon;
   Packet pkt;
   driver drv;
   //DUT
   RamChip #(4,8)DUT(iftest.Address, iftest.Data, iftest.CS, iftest.WE, iftest.OE);

   initial clk=0;

   always #5 clk = ~clk;

   initial begin
      mon = new();
      drv = new(iftest);
      repeat(8) begin
	 pkt = new();
	 assert(pkt.randomize());
	 drv.send_rqt(pkt);
      end
   end
   
   

endmodule // top




































