// Code your testbench here
// or browse Examples

import uvm_pkg::*;
`include "uvm_macros.svh"


`include "test.sv"


