// Code your testbench here
// or browse Examples


import uvm_pkg::*;
`include "uvm_macros.svh"

`include "mem.v"
`include "read_if.sv"
`include "write_if.sv"

`include "top.sv"
`include "rw_seq_item.sv"
`include "rw_sequence.sv"
`include "v_sequencer.sv"
`include "rw_driver.sv"
`include "rw_agent.sv"
`include "rw_env.sv"
`include "rw_test.sv"