abhaysingh@Abhays-MacBook-Pro.local.8994