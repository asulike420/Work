// Code your testbench here
// or browse Examples


`include "reg_defs.sv"
`include "ahb_if.sv"
`include "mem_ss.sv"
`include "mem_ss_wrapper.sv"
`include "ahb_agent_pkg.sv"
`include "mem_ss_reg_pkg.sv"


`include "mem_ss_env_pkg.sv"

`include "mem_ss_seq_lib_pkg.sv"
`include "mem_ss_test_lib_pkg.sv"
`include "top_tb.sv"