package router_stimulus_pkg;

import uvm_pkg::*;

`include "packet.sv"

// Lab 2: Task 7, Step 2 - include the packet_sequence.sv file
//
// ToDo



// Lab 2: Task 9, Step 2 - include the packet_da_3.sv file
//
// ToDo



endpackage
