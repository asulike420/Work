// Code your design here
`include "host_io.sv"
`include "router_io.sv"
`include "reset_io.sv"
`include "router.sv"
`include "router_test_top.sv"

