
1. Port coresponding to Data received from 2 channels
2. Port coresponding  Output captured from 1 channel
3. Common queue to track the order in wich data is captured  from the input channels
  Item in the queue must contain the data and the timestamp
4. Expected queue


  1. continius stream of data in both the channels
    a) starting at the same time
    b) starting at different times

  2. arbitary data
   

  
    
 
